`ifndef UART_COMM_
`define UART_COMM_
//`timescale 1ns / 1ps
`include "buffer.v"
//`include "fifo.v"
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/06/15 07:07:54
// Design Name: 
// Module Name: uart_comm
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module uart_comm 
	#(
    parameter ID = 1,
	parameter BAUDRATE = 9600,
	parameter CLOCKRATE = 100000000
	)(
	input CLK,
	input RST,
	
	input send_flag,
	input [7:0] send_data,
	input recv_flag,
	output [7:0] recv_data,

    output send_ack, recv_ack,
    //output reg send_ack, recv_ack,
	output sendable,
	output receivable,
	
	output reg Tx,
	input Rx
    );

	reg recv_write_flag;
	reg [7:0] recv_write_data;
	wire recv_empty, recv_full, rbuf_rack, rbuf_wack, rbuf_a;
	//fifo #(.WIDTH(8)) recv_buffer(CLK, RST, recv_flag, recv_data, recv_write_flag, recv_write_data, recv_empty, recv_full);
    buffer#(.BUF_ID(ID+10),.ADDR_L(5),.DATA_L(8)) recv_buffer
    (CLK,RST,recv_flag,recv_write_flag,recv_write_data,recv_data,/*rbuf_rack*/recv_ack,rbuf_wack,rbuf_a,recv_full);
    assign recv_empty = ~rbuf_a;
	reg send_read_flag;
	wire [7:0] send_read_data;
	reg [7:0] send_read_data_buf;
	wire send_empty, send_full, sbuf_rack, sbuf_wack, sbuf_a;
	//fifo #(.WIDTH(8)) send_buffer(CLK, RST, send_read_flag, send_read_data, send_flag, send_data, send_empty, send_full);
    buffer#(.BUF_ID(ID+11),.ADDR_L(5),.DATA_L(8)) send_buffer
    (CLK,RST,send_read_flag,send_flag,send_data,send_read_data,sbuf_rack,/*sbuf_wack*/send_ack,sbuf_a,send_full);
    assign send_empty = ~sbuf_a;
	//assign receivable = !recv_empty;
	assign receivable = rbuf_a;
	assign sendable = !send_full;
	
	localparam SAMPLE_INTERVAL = CLOCKRATE / BAUDRATE;
	
	localparam STATUS_IDLE = 0;
	localparam STATUS_BEGIN = 1;
	localparam STATUS_DATA = 2;
	localparam STATUS_VALID = 4;
	localparam STATUS_END = 8;
	reg [3:0] recv_status;
	reg [2:0] recv_bit;
	reg recv_parity;
	
	integer recv_counter;
	reg recv_clock;
	
	wire sample = recv_counter == SAMPLE_INTERVAL / 2;
	
	always @(posedge CLK or posedge RST) begin
		if(RST) begin
			recv_write_flag <= 0;
			recv_write_data <= 0;
			recv_status <= STATUS_IDLE;
			recv_bit <= 0;
			recv_parity <= 0;
			recv_counter <= 0;
			recv_clock <= 0;
            //recv_ack = 0;
		end else begin
            //recv_ack = 0;
			//recv_write_flag <= 0;
			if(recv_clock) begin
				if(recv_counter == SAMPLE_INTERVAL - 1)
					recv_counter <= 0;
				else
					recv_counter <= recv_counter + 1;
			end
			if(recv_status == STATUS_IDLE) begin
				if(!Rx) begin
					recv_status <= STATUS_BEGIN;
					recv_counter <= 0;
					recv_clock <= 1;
				end
			end else if(sample) begin
				case(recv_status)
				STATUS_BEGIN:begin
					if(!Rx) begin
						recv_status <= STATUS_DATA;
						recv_bit <= 0;
						recv_parity <= 0;
					end else begin
						recv_status <= STATUS_IDLE;
						recv_clock <= 0;
					end
				end
				
				STATUS_DATA:begin
                    //$display("UART:%0d Recv bit %b",ID,Rx);
					recv_parity <= recv_parity ^ Rx;
					recv_write_data[recv_bit] <= Rx;
					recv_bit <= recv_bit + 1;
					if(recv_bit == 7)
						recv_status <= STATUS_VALID;
				end
				
				STATUS_VALID:begin
					if(recv_parity == Rx && !recv_full)
						recv_write_flag <= 1;
					recv_status <= STATUS_END;
				end
				
				STATUS_END: begin
                    //$display("UART:%0d Received %b",ID,recv_write_data);
					recv_status <= STATUS_IDLE;
					recv_clock <= 0;
                    //recv_ack = 1;
				end
				endcase
			end
		end
	end

    always @(posedge rbuf_wack) begin
        recv_write_flag <= 0;
    end
	
	integer counter;
	always @(posedge CLK or posedge RST) begin
		if(RST) begin
			counter <= 0;
		end else begin
			counter <= counter + 1;
			if(counter == SAMPLE_INTERVAL - 1)
				counter <= 0;
		end
	end
	
	reg [3:0] send_status;
	reg [2:0] send_bit;
	reg send_parity;
	reg tosend;
	
	always @(posedge CLK or posedge RST) begin
		if(RST) begin
			send_read_flag <= 0;
			send_read_data_buf <= 0;
			send_status <= STATUS_IDLE;
			send_bit <= 0;
			send_parity <= 0;
			tosend <= 0;
			Tx <= 1;
            //send_ack = 0;
		end else begin
			//send_read_flag <= 0;
			//send_ack = 0;	
			if(counter == 0) begin
				case(send_status)
				STATUS_IDLE:begin
					//if(!send_empty) begin
					if(sbuf_a) begin
						//send_read_data_buf <= send_read_data;
						send_read_flag = 1;
						Tx <= 0;
						//send_status <= STATUS_DATA;
						send_bit <= 0;
						send_parity <= 0;
					end
				end
				
				STATUS_DATA:begin
                    //$display("UART:%0d Send bit %b",ID,send_read_data_buf[send_bit]);
					Tx <= send_read_data_buf[send_bit];
					send_parity <= send_parity ^ send_read_data_buf[send_bit];
					send_bit <= send_bit + 1;
					if(send_bit == 7)
						send_status <= STATUS_VALID;
				end
				
				STATUS_VALID:begin
					Tx <= send_parity;
					send_status <= STATUS_END;
				end
				
				STATUS_END:begin
                    //$display("UART:%0d Sent %b",ID,send_read_data_buf);
                    //send_ack = 1;
					Tx <= 1;
					send_status <= STATUS_IDLE;
					tosend = 0;
				end
				endcase
			end
		end
	end

    always @(posedge sbuf_rack) begin
        send_status <= STATUS_DATA;
		send_read_data_buf <= send_read_data;
        send_read_flag <= 0;
    end

endmodule
`endif
